
module niosLab2 (
	clk_clk,
	leds_name,
	reset_reset_n,
	fases_phases);	

	input		clk_clk;
	output	[3:0]	leds_name;
	input		reset_reset_n;
	output	[3:0]	fases_phases;
endmodule
