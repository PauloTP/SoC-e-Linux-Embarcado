-- niosLab2_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosLab2_tb is
end entity niosLab2_tb;

architecture rtl of niosLab2_tb is
	component niosLab2 is
		port (
			clk_clk         : in  std_logic                    := 'X';             -- clk
			leds_name       : out std_logic_vector(3 downto 0);                    -- name
			reset_reset_n   : in  std_logic                    := 'X';             -- reset_n
			switches_export : in  std_logic_vector(5 downto 0) := (others => 'X')  -- export
		);
	end component niosLab2;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			clk      : in std_logic                    := 'X';             -- clk
			sig_name : in std_logic_vector(3 downto 0) := (others => 'X'); -- name
			reset    : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : out std_logic_vector(5 downto 0)   -- export
		);
	end component altera_conduit_bfm_0002;

	signal nioslab2_inst_clk_bfm_clk_clk             : std_logic;                    -- niosLab2_inst_clk_bfm:clk -> [niosLab2_inst:clk_clk, niosLab2_inst_leds_bfm:clk, niosLab2_inst_reset_bfm:clk]
	signal nioslab2_inst_leds_name                   : std_logic_vector(3 downto 0); -- niosLab2_inst:leds_name -> niosLab2_inst_leds_bfm:sig_name
	signal nioslab2_inst_switches_bfm_conduit_export : std_logic_vector(5 downto 0); -- niosLab2_inst_switches_bfm:sig_export -> niosLab2_inst:switches_export
	signal nioslab2_inst_reset_bfm_reset_reset       : std_logic;                    -- niosLab2_inst_reset_bfm:reset -> niosLab2_inst:reset_reset_n

begin

	nioslab2_inst : component niosLab2
		port map (
			clk_clk         => nioslab2_inst_clk_bfm_clk_clk,             --      clk.clk
			leds_name       => nioslab2_inst_leds_name,                   --     leds.name
			reset_reset_n   => nioslab2_inst_reset_bfm_reset_reset,       --    reset.reset_n
			switches_export => nioslab2_inst_switches_bfm_conduit_export  -- switches.export
		);

	nioslab2_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nioslab2_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nioslab2_inst_leds_bfm : component altera_conduit_bfm
		port map (
			clk      => nioslab2_inst_clk_bfm_clk_clk, --     clk.clk
			sig_name => nioslab2_inst_leds_name,       -- conduit.name
			reset    => '0'                            -- (terminated)
		);

	nioslab2_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nioslab2_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => nioslab2_inst_clk_bfm_clk_clk        --   clk.clk
		);

	nioslab2_inst_switches_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nioslab2_inst_switches_bfm_conduit_export  -- conduit.export
		);

end architecture rtl; -- of niosLab2_tb
